magic
tech sky130A
timestamp 1743271696
<< pwell >>
rect -692 -150 692 150
<< nnmos >>
rect -578 -21 -528 21
rect -499 -21 -449 21
rect -420 -21 -370 21
rect -341 -21 -291 21
rect -262 -21 -212 21
rect -183 -21 -133 21
rect -104 -21 -54 21
rect -25 -21 25 21
rect 54 -21 104 21
rect 133 -21 183 21
rect 212 -21 262 21
rect 291 -21 341 21
rect 370 -21 420 21
rect 449 -21 499 21
rect 528 -21 578 21
<< mvndiff >>
rect -607 15 -578 21
rect -607 -15 -601 15
rect -584 -15 -578 15
rect -607 -21 -578 -15
rect -528 15 -499 21
rect -528 -15 -522 15
rect -505 -15 -499 15
rect -528 -21 -499 -15
rect -449 15 -420 21
rect -449 -15 -443 15
rect -426 -15 -420 15
rect -449 -21 -420 -15
rect -370 15 -341 21
rect -370 -15 -364 15
rect -347 -15 -341 15
rect -370 -21 -341 -15
rect -291 15 -262 21
rect -291 -15 -285 15
rect -268 -15 -262 15
rect -291 -21 -262 -15
rect -212 15 -183 21
rect -212 -15 -206 15
rect -189 -15 -183 15
rect -212 -21 -183 -15
rect -133 15 -104 21
rect -133 -15 -127 15
rect -110 -15 -104 15
rect -133 -21 -104 -15
rect -54 15 -25 21
rect -54 -15 -48 15
rect -31 -15 -25 15
rect -54 -21 -25 -15
rect 25 15 54 21
rect 25 -15 31 15
rect 48 -15 54 15
rect 25 -21 54 -15
rect 104 15 133 21
rect 104 -15 110 15
rect 127 -15 133 15
rect 104 -21 133 -15
rect 183 15 212 21
rect 183 -15 189 15
rect 206 -15 212 15
rect 183 -21 212 -15
rect 262 15 291 21
rect 262 -15 268 15
rect 285 -15 291 15
rect 262 -21 291 -15
rect 341 15 370 21
rect 341 -15 347 15
rect 364 -15 370 15
rect 341 -21 370 -15
rect 420 15 449 21
rect 420 -15 426 15
rect 443 -15 449 15
rect 420 -21 449 -15
rect 499 15 528 21
rect 499 -15 505 15
rect 522 -15 528 15
rect 499 -21 528 -15
rect 578 15 607 21
rect 578 -15 584 15
rect 601 -15 607 15
rect 578 -21 607 -15
<< mvndiffc >>
rect -601 -15 -584 15
rect -522 -15 -505 15
rect -443 -15 -426 15
rect -364 -15 -347 15
rect -285 -15 -268 15
rect -206 -15 -189 15
rect -127 -15 -110 15
rect -48 -15 -31 15
rect 31 -15 48 15
rect 110 -15 127 15
rect 189 -15 206 15
rect 268 -15 285 15
rect 347 -15 364 15
rect 426 -15 443 15
rect 505 -15 522 15
rect 584 -15 601 15
<< mvpsubdiff >>
rect -674 126 674 132
rect -674 109 -620 126
rect 620 109 674 126
rect -674 103 674 109
rect -674 78 -645 103
rect -674 -78 -668 78
rect -651 -78 -645 78
rect 645 78 674 103
rect -674 -103 -645 -78
rect 645 -78 651 78
rect 668 -78 674 78
rect 645 -103 674 -78
rect -674 -109 674 -103
rect -674 -126 -620 -109
rect 620 -126 674 -109
rect -674 -132 674 -126
<< mvpsubdiffcont >>
rect -620 109 620 126
rect -668 -78 -651 78
rect 651 -78 668 78
rect -620 -126 620 -109
<< poly >>
rect -578 57 -528 65
rect -578 40 -570 57
rect -536 40 -528 57
rect -578 21 -528 40
rect -499 57 -449 65
rect -499 40 -491 57
rect -457 40 -449 57
rect -499 21 -449 40
rect -420 57 -370 65
rect -420 40 -412 57
rect -378 40 -370 57
rect -420 21 -370 40
rect -341 57 -291 65
rect -341 40 -333 57
rect -299 40 -291 57
rect -341 21 -291 40
rect -262 57 -212 65
rect -262 40 -254 57
rect -220 40 -212 57
rect -262 21 -212 40
rect -183 57 -133 65
rect -183 40 -175 57
rect -141 40 -133 57
rect -183 21 -133 40
rect -104 57 -54 65
rect -104 40 -96 57
rect -62 40 -54 57
rect -104 21 -54 40
rect -25 57 25 65
rect -25 40 -17 57
rect 17 40 25 57
rect -25 21 25 40
rect 54 57 104 65
rect 54 40 62 57
rect 96 40 104 57
rect 54 21 104 40
rect 133 57 183 65
rect 133 40 141 57
rect 175 40 183 57
rect 133 21 183 40
rect 212 57 262 65
rect 212 40 220 57
rect 254 40 262 57
rect 212 21 262 40
rect 291 57 341 65
rect 291 40 299 57
rect 333 40 341 57
rect 291 21 341 40
rect 370 57 420 65
rect 370 40 378 57
rect 412 40 420 57
rect 370 21 420 40
rect 449 57 499 65
rect 449 40 457 57
rect 491 40 499 57
rect 449 21 499 40
rect 528 57 578 65
rect 528 40 536 57
rect 570 40 578 57
rect 528 21 578 40
rect -578 -40 -528 -21
rect -578 -57 -570 -40
rect -536 -57 -528 -40
rect -578 -65 -528 -57
rect -499 -40 -449 -21
rect -499 -57 -491 -40
rect -457 -57 -449 -40
rect -499 -65 -449 -57
rect -420 -40 -370 -21
rect -420 -57 -412 -40
rect -378 -57 -370 -40
rect -420 -65 -370 -57
rect -341 -40 -291 -21
rect -341 -57 -333 -40
rect -299 -57 -291 -40
rect -341 -65 -291 -57
rect -262 -40 -212 -21
rect -262 -57 -254 -40
rect -220 -57 -212 -40
rect -262 -65 -212 -57
rect -183 -40 -133 -21
rect -183 -57 -175 -40
rect -141 -57 -133 -40
rect -183 -65 -133 -57
rect -104 -40 -54 -21
rect -104 -57 -96 -40
rect -62 -57 -54 -40
rect -104 -65 -54 -57
rect -25 -40 25 -21
rect -25 -57 -17 -40
rect 17 -57 25 -40
rect -25 -65 25 -57
rect 54 -40 104 -21
rect 54 -57 62 -40
rect 96 -57 104 -40
rect 54 -65 104 -57
rect 133 -40 183 -21
rect 133 -57 141 -40
rect 175 -57 183 -40
rect 133 -65 183 -57
rect 212 -40 262 -21
rect 212 -57 220 -40
rect 254 -57 262 -40
rect 212 -65 262 -57
rect 291 -40 341 -21
rect 291 -57 299 -40
rect 333 -57 341 -40
rect 291 -65 341 -57
rect 370 -40 420 -21
rect 370 -57 378 -40
rect 412 -57 420 -40
rect 370 -65 420 -57
rect 449 -40 499 -21
rect 449 -57 457 -40
rect 491 -57 499 -40
rect 449 -65 499 -57
rect 528 -40 578 -21
rect 528 -57 536 -40
rect 570 -57 578 -40
rect 528 -65 578 -57
<< polycont >>
rect -570 40 -536 57
rect -491 40 -457 57
rect -412 40 -378 57
rect -333 40 -299 57
rect -254 40 -220 57
rect -175 40 -141 57
rect -96 40 -62 57
rect -17 40 17 57
rect 62 40 96 57
rect 141 40 175 57
rect 220 40 254 57
rect 299 40 333 57
rect 378 40 412 57
rect 457 40 491 57
rect 536 40 570 57
rect -570 -57 -536 -40
rect -491 -57 -457 -40
rect -412 -57 -378 -40
rect -333 -57 -299 -40
rect -254 -57 -220 -40
rect -175 -57 -141 -40
rect -96 -57 -62 -40
rect -17 -57 17 -40
rect 62 -57 96 -40
rect 141 -57 175 -40
rect 220 -57 254 -40
rect 299 -57 333 -40
rect 378 -57 412 -40
rect 457 -57 491 -40
rect 536 -57 570 -40
<< locali >>
rect -668 109 -620 126
rect 620 109 668 126
rect -668 78 -651 109
rect 651 78 668 109
rect -578 40 -570 57
rect -536 40 -528 57
rect -499 40 -491 57
rect -457 40 -449 57
rect -420 40 -412 57
rect -378 40 -370 57
rect -341 40 -333 57
rect -299 40 -291 57
rect -262 40 -254 57
rect -220 40 -212 57
rect -183 40 -175 57
rect -141 40 -133 57
rect -104 40 -96 57
rect -62 40 -54 57
rect -25 40 -17 57
rect 17 40 25 57
rect 54 40 62 57
rect 96 40 104 57
rect 133 40 141 57
rect 175 40 183 57
rect 212 40 220 57
rect 254 40 262 57
rect 291 40 299 57
rect 333 40 341 57
rect 370 40 378 57
rect 412 40 420 57
rect 449 40 457 57
rect 491 40 499 57
rect 528 40 536 57
rect 570 40 578 57
rect -601 15 -584 23
rect -601 -23 -584 -15
rect -522 15 -505 23
rect -522 -23 -505 -15
rect -443 15 -426 23
rect -443 -23 -426 -15
rect -364 15 -347 23
rect -364 -23 -347 -15
rect -285 15 -268 23
rect -285 -23 -268 -15
rect -206 15 -189 23
rect -206 -23 -189 -15
rect -127 15 -110 23
rect -127 -23 -110 -15
rect -48 15 -31 23
rect -48 -23 -31 -15
rect 31 15 48 23
rect 31 -23 48 -15
rect 110 15 127 23
rect 110 -23 127 -15
rect 189 15 206 23
rect 189 -23 206 -15
rect 268 15 285 23
rect 268 -23 285 -15
rect 347 15 364 23
rect 347 -23 364 -15
rect 426 15 443 23
rect 426 -23 443 -15
rect 505 15 522 23
rect 505 -23 522 -15
rect 584 15 601 23
rect 584 -23 601 -15
rect -578 -57 -570 -40
rect -536 -57 -528 -40
rect -499 -57 -491 -40
rect -457 -57 -449 -40
rect -420 -57 -412 -40
rect -378 -57 -370 -40
rect -341 -57 -333 -40
rect -299 -57 -291 -40
rect -262 -57 -254 -40
rect -220 -57 -212 -40
rect -183 -57 -175 -40
rect -141 -57 -133 -40
rect -104 -57 -96 -40
rect -62 -57 -54 -40
rect -25 -57 -17 -40
rect 17 -57 25 -40
rect 54 -57 62 -40
rect 96 -57 104 -40
rect 133 -57 141 -40
rect 175 -57 183 -40
rect 212 -57 220 -40
rect 254 -57 262 -40
rect 291 -57 299 -40
rect 333 -57 341 -40
rect 370 -57 378 -40
rect 412 -57 420 -40
rect 449 -57 457 -40
rect 491 -57 499 -40
rect 528 -57 536 -40
rect 570 -57 578 -40
rect -668 -109 -651 -78
rect 651 -109 668 -78
rect -668 -126 -620 -109
rect 620 -126 668 -109
<< viali >>
rect -570 40 -536 57
rect -491 40 -457 57
rect -412 40 -378 57
rect -333 40 -299 57
rect -254 40 -220 57
rect -175 40 -141 57
rect -96 40 -62 57
rect -17 40 17 57
rect 62 40 96 57
rect 141 40 175 57
rect 220 40 254 57
rect 299 40 333 57
rect 378 40 412 57
rect 457 40 491 57
rect 536 40 570 57
rect -601 -15 -584 15
rect -522 -15 -505 15
rect -443 -15 -426 15
rect -364 -15 -347 15
rect -285 -15 -268 15
rect -206 -15 -189 15
rect -127 -15 -110 15
rect -48 -15 -31 15
rect 31 -15 48 15
rect 110 -15 127 15
rect 189 -15 206 15
rect 268 -15 285 15
rect 347 -15 364 15
rect 426 -15 443 15
rect 505 -15 522 15
rect 584 -15 601 15
rect -570 -57 -536 -40
rect -491 -57 -457 -40
rect -412 -57 -378 -40
rect -333 -57 -299 -40
rect -254 -57 -220 -40
rect -175 -57 -141 -40
rect -96 -57 -62 -40
rect -17 -57 17 -40
rect 62 -57 96 -40
rect 141 -57 175 -40
rect 220 -57 254 -40
rect 299 -57 333 -40
rect 378 -57 412 -40
rect 457 -57 491 -40
rect 536 -57 570 -40
<< metal1 >>
rect -576 57 -530 60
rect -576 40 -570 57
rect -536 40 -530 57
rect -576 37 -530 40
rect -497 57 -451 60
rect -497 40 -491 57
rect -457 40 -451 57
rect -497 37 -451 40
rect -418 57 -372 60
rect -418 40 -412 57
rect -378 40 -372 57
rect -418 37 -372 40
rect -339 57 -293 60
rect -339 40 -333 57
rect -299 40 -293 57
rect -339 37 -293 40
rect -260 57 -214 60
rect -260 40 -254 57
rect -220 40 -214 57
rect -260 37 -214 40
rect -181 57 -135 60
rect -181 40 -175 57
rect -141 40 -135 57
rect -181 37 -135 40
rect -102 57 -56 60
rect -102 40 -96 57
rect -62 40 -56 57
rect -102 37 -56 40
rect -23 57 23 60
rect -23 40 -17 57
rect 17 40 23 57
rect -23 37 23 40
rect 56 57 102 60
rect 56 40 62 57
rect 96 40 102 57
rect 56 37 102 40
rect 135 57 181 60
rect 135 40 141 57
rect 175 40 181 57
rect 135 37 181 40
rect 214 57 260 60
rect 214 40 220 57
rect 254 40 260 57
rect 214 37 260 40
rect 293 57 339 60
rect 293 40 299 57
rect 333 40 339 57
rect 293 37 339 40
rect 372 57 418 60
rect 372 40 378 57
rect 412 40 418 57
rect 372 37 418 40
rect 451 57 497 60
rect 451 40 457 57
rect 491 40 497 57
rect 451 37 497 40
rect 530 57 576 60
rect 530 40 536 57
rect 570 40 576 57
rect 530 37 576 40
rect -604 15 -581 21
rect -604 -15 -601 15
rect -584 -15 -581 15
rect -604 -21 -581 -15
rect -525 15 -502 21
rect -525 -15 -522 15
rect -505 -15 -502 15
rect -525 -21 -502 -15
rect -446 15 -423 21
rect -446 -15 -443 15
rect -426 -15 -423 15
rect -446 -21 -423 -15
rect -367 15 -344 21
rect -367 -15 -364 15
rect -347 -15 -344 15
rect -367 -21 -344 -15
rect -288 15 -265 21
rect -288 -15 -285 15
rect -268 -15 -265 15
rect -288 -21 -265 -15
rect -209 15 -186 21
rect -209 -15 -206 15
rect -189 -15 -186 15
rect -209 -21 -186 -15
rect -130 15 -107 21
rect -130 -15 -127 15
rect -110 -15 -107 15
rect -130 -21 -107 -15
rect -51 15 -28 21
rect -51 -15 -48 15
rect -31 -15 -28 15
rect -51 -21 -28 -15
rect 28 15 51 21
rect 28 -15 31 15
rect 48 -15 51 15
rect 28 -21 51 -15
rect 107 15 130 21
rect 107 -15 110 15
rect 127 -15 130 15
rect 107 -21 130 -15
rect 186 15 209 21
rect 186 -15 189 15
rect 206 -15 209 15
rect 186 -21 209 -15
rect 265 15 288 21
rect 265 -15 268 15
rect 285 -15 288 15
rect 265 -21 288 -15
rect 344 15 367 21
rect 344 -15 347 15
rect 364 -15 367 15
rect 344 -21 367 -15
rect 423 15 446 21
rect 423 -15 426 15
rect 443 -15 446 15
rect 423 -21 446 -15
rect 502 15 525 21
rect 502 -15 505 15
rect 522 -15 525 15
rect 502 -21 525 -15
rect 581 15 604 21
rect 581 -15 584 15
rect 601 -15 604 15
rect 581 -21 604 -15
rect -576 -40 -530 -37
rect -576 -57 -570 -40
rect -536 -57 -530 -40
rect -576 -60 -530 -57
rect -497 -40 -451 -37
rect -497 -57 -491 -40
rect -457 -57 -451 -40
rect -497 -60 -451 -57
rect -418 -40 -372 -37
rect -418 -57 -412 -40
rect -378 -57 -372 -40
rect -418 -60 -372 -57
rect -339 -40 -293 -37
rect -339 -57 -333 -40
rect -299 -57 -293 -40
rect -339 -60 -293 -57
rect -260 -40 -214 -37
rect -260 -57 -254 -40
rect -220 -57 -214 -40
rect -260 -60 -214 -57
rect -181 -40 -135 -37
rect -181 -57 -175 -40
rect -141 -57 -135 -40
rect -181 -60 -135 -57
rect -102 -40 -56 -37
rect -102 -57 -96 -40
rect -62 -57 -56 -40
rect -102 -60 -56 -57
rect -23 -40 23 -37
rect -23 -57 -17 -40
rect 17 -57 23 -40
rect -23 -60 23 -57
rect 56 -40 102 -37
rect 56 -57 62 -40
rect 96 -57 102 -40
rect 56 -60 102 -57
rect 135 -40 181 -37
rect 135 -57 141 -40
rect 175 -57 181 -40
rect 135 -60 181 -57
rect 214 -40 260 -37
rect 214 -57 220 -40
rect 254 -57 260 -40
rect 214 -60 260 -57
rect 293 -40 339 -37
rect 293 -57 299 -40
rect 333 -57 339 -40
rect 293 -60 339 -57
rect 372 -40 418 -37
rect 372 -57 378 -40
rect 412 -57 418 -40
rect 372 -60 418 -57
rect 451 -40 497 -37
rect 451 -57 457 -40
rect 491 -57 497 -40
rect 451 -60 497 -57
rect 530 -40 576 -37
rect 530 -57 536 -40
rect 570 -57 576 -40
rect 530 -60 576 -57
<< properties >>
string FIXED_BBOX -659 -117 659 117
string gencell sky130_fd_pr__nfet_03v3_nvt
string library sky130
string parameters w 0.420 l 0.50 m 1 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
