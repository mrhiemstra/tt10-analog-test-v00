MACRO sky130_fd_pr__nfet_03v3_nvt_PDAVVX
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__nfet_03v3_nvt_PDAVVX ;
  ORIGIN 6.595 1.175 ;
  SIZE 13.190 BY 2.350 ;
  OBS
      LAYER pwell ;
        RECT -6.920 -1.500 6.920 1.500 ;
      LAYER li1 ;
        RECT -6.680 1.090 6.680 1.260 ;
        RECT -6.680 -1.090 -6.510 1.090 ;
        RECT -5.780 0.400 -5.280 0.570 ;
        RECT -4.990 0.400 -4.490 0.570 ;
        RECT -4.200 0.400 -3.700 0.570 ;
        RECT -3.410 0.400 -2.910 0.570 ;
        RECT -2.620 0.400 -2.120 0.570 ;
        RECT -1.830 0.400 -1.330 0.570 ;
        RECT -1.040 0.400 -0.540 0.570 ;
        RECT -0.250 0.400 0.250 0.570 ;
        RECT 0.540 0.400 1.040 0.570 ;
        RECT 1.330 0.400 1.830 0.570 ;
        RECT 2.120 0.400 2.620 0.570 ;
        RECT 2.910 0.400 3.410 0.570 ;
        RECT 3.700 0.400 4.200 0.570 ;
        RECT 4.490 0.400 4.990 0.570 ;
        RECT 5.280 0.400 5.780 0.570 ;
        RECT -6.010 -0.230 -5.840 0.230 ;
        RECT -5.220 -0.230 -5.050 0.230 ;
        RECT -4.430 -0.230 -4.260 0.230 ;
        RECT -3.640 -0.230 -3.470 0.230 ;
        RECT -2.850 -0.230 -2.680 0.230 ;
        RECT -2.060 -0.230 -1.890 0.230 ;
        RECT -1.270 -0.230 -1.100 0.230 ;
        RECT -0.480 -0.230 -0.310 0.230 ;
        RECT 0.310 -0.230 0.480 0.230 ;
        RECT 1.100 -0.230 1.270 0.230 ;
        RECT 1.890 -0.230 2.060 0.230 ;
        RECT 2.680 -0.230 2.850 0.230 ;
        RECT 3.470 -0.230 3.640 0.230 ;
        RECT 4.260 -0.230 4.430 0.230 ;
        RECT 5.050 -0.230 5.220 0.230 ;
        RECT 5.840 -0.230 6.010 0.230 ;
        RECT -5.780 -0.570 -5.280 -0.400 ;
        RECT -4.990 -0.570 -4.490 -0.400 ;
        RECT -4.200 -0.570 -3.700 -0.400 ;
        RECT -3.410 -0.570 -2.910 -0.400 ;
        RECT -2.620 -0.570 -2.120 -0.400 ;
        RECT -1.830 -0.570 -1.330 -0.400 ;
        RECT -1.040 -0.570 -0.540 -0.400 ;
        RECT -0.250 -0.570 0.250 -0.400 ;
        RECT 0.540 -0.570 1.040 -0.400 ;
        RECT 1.330 -0.570 1.830 -0.400 ;
        RECT 2.120 -0.570 2.620 -0.400 ;
        RECT 2.910 -0.570 3.410 -0.400 ;
        RECT 3.700 -0.570 4.200 -0.400 ;
        RECT 4.490 -0.570 4.990 -0.400 ;
        RECT 5.280 -0.570 5.780 -0.400 ;
        RECT 6.510 -1.090 6.680 1.090 ;
        RECT -6.680 -1.260 6.680 -1.090 ;
      LAYER met1 ;
        RECT -5.760 0.370 -5.300 0.600 ;
        RECT -4.970 0.370 -4.510 0.600 ;
        RECT -4.180 0.370 -3.720 0.600 ;
        RECT -3.390 0.370 -2.930 0.600 ;
        RECT -2.600 0.370 -2.140 0.600 ;
        RECT -1.810 0.370 -1.350 0.600 ;
        RECT -1.020 0.370 -0.560 0.600 ;
        RECT -0.230 0.370 0.230 0.600 ;
        RECT 0.560 0.370 1.020 0.600 ;
        RECT 1.350 0.370 1.810 0.600 ;
        RECT 2.140 0.370 2.600 0.600 ;
        RECT 2.930 0.370 3.390 0.600 ;
        RECT 3.720 0.370 4.180 0.600 ;
        RECT 4.510 0.370 4.970 0.600 ;
        RECT 5.300 0.370 5.760 0.600 ;
        RECT -6.040 -0.210 -5.810 0.210 ;
        RECT -5.250 -0.210 -5.020 0.210 ;
        RECT -4.460 -0.210 -4.230 0.210 ;
        RECT -3.670 -0.210 -3.440 0.210 ;
        RECT -2.880 -0.210 -2.650 0.210 ;
        RECT -2.090 -0.210 -1.860 0.210 ;
        RECT -1.300 -0.210 -1.070 0.210 ;
        RECT -0.510 -0.210 -0.280 0.210 ;
        RECT 0.280 -0.210 0.510 0.210 ;
        RECT 1.070 -0.210 1.300 0.210 ;
        RECT 1.860 -0.210 2.090 0.210 ;
        RECT 2.650 -0.210 2.880 0.210 ;
        RECT 3.440 -0.210 3.670 0.210 ;
        RECT 4.230 -0.210 4.460 0.210 ;
        RECT 5.020 -0.210 5.250 0.210 ;
        RECT 5.810 -0.210 6.040 0.210 ;
        RECT -5.760 -0.600 -5.300 -0.370 ;
        RECT -4.970 -0.600 -4.510 -0.370 ;
        RECT -4.180 -0.600 -3.720 -0.370 ;
        RECT -3.390 -0.600 -2.930 -0.370 ;
        RECT -2.600 -0.600 -2.140 -0.370 ;
        RECT -1.810 -0.600 -1.350 -0.370 ;
        RECT -1.020 -0.600 -0.560 -0.370 ;
        RECT -0.230 -0.600 0.230 -0.370 ;
        RECT 0.560 -0.600 1.020 -0.370 ;
        RECT 1.350 -0.600 1.810 -0.370 ;
        RECT 2.140 -0.600 2.600 -0.370 ;
        RECT 2.930 -0.600 3.390 -0.370 ;
        RECT 3.720 -0.600 4.180 -0.370 ;
        RECT 4.510 -0.600 4.970 -0.370 ;
        RECT 5.300 -0.600 5.760 -0.370 ;
  END
END sky130_fd_pr__nfet_03v3_nvt_PDAVVX
END LIBRARY

